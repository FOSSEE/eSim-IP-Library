module xor21(c,a,b);
input a,b;
output c;
xor (c,a,b);
endmodule
